-- Memory.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Memory is
	port (
		clk_clk            : in  std_logic                     := '0';             --    clk.clk
		reset_reset        : in  std_logic                     := '0';             --  reset.reset
		reset_reset_req    : in  std_logic                     := '0';             --       .reset_req
		sortie_address     : in  std_logic_vector(7 downto 0)  := (others => '0'); -- sortie.address
		sortie_debugaccess : in  std_logic                     := '0';             --       .debugaccess
		sortie_clken       : in  std_logic                     := '0';             --       .clken
		sortie_chipselect  : in  std_logic                     := '0';             --       .chipselect
		sortie_write       : in  std_logic                     := '0';             --       .write
		sortie_readdata    : out std_logic_vector(15 downto 0);                    --       .readdata
		sortie_writedata   : in  std_logic_vector(15 downto 0) := (others => '0'); --       .writedata
		sortie_byteenable  : in  std_logic_vector(1 downto 0)  := (others => '0')  --       .byteenable
	);
end entity Memory;

architecture rtl of Memory is
	component Memory_onchip_memory2_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			debugaccess : in  std_logic                     := 'X';             -- debugaccess
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(15 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component Memory_onchip_memory2_0;

begin

	onchip_memory2_0 : component Memory_onchip_memory2_0
		port map (
			clk         => clk_clk,            --   clk1.clk
			address     => sortie_address,     --     s1.address
			debugaccess => sortie_debugaccess, --       .debugaccess
			clken       => sortie_clken,       --       .clken
			chipselect  => sortie_chipselect,  --       .chipselect
			write       => sortie_write,       --       .write
			readdata    => sortie_readdata,    --       .readdata
			writedata   => sortie_writedata,   --       .writedata
			byteenable  => sortie_byteenable,  --       .byteenable
			reset       => reset_reset,        -- reset1.reset
			reset_req   => reset_reset_req     --       .reset_req
		);

end architecture rtl; -- of Memory
